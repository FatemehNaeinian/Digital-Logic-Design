`timescale 1ns/1ns
module NAND_GATE_TESTBENCH();
  logic aa=1; 
  logic bb=1;
  wire ww;
  NAND_GATE UUT(aa,bb,ww);
  initial begin
  #20 aa=0;
  #20 aa=1;
  #20 bb=0;
  #20 bb=1;
  #20 aa=0 ;bb=0;
  #20 aa=1 ;bb=0;
  #20   $stop;
  end 
endmodule