`timescale 1ns/1ns
module barrel16 (input [15:0]M,[3:0]S , output SHO[15:0]);
mux16to1 T1({M[0],M[1],M[2],M[3],M[4],M[5],M[6],M[7],M[8],M[9],M[10],M[11],M[12],M[13],M[14],M[15]},S,SHO[0]);
mux16to1 T2({M[1],M[2],M[3],M[4],M[5],M[6],M[7],M[8],M[9],M[10],M[11],M[12],M[13],M[14],M[15],M[0]},S,SHO[1]);
mux16to1 T3({M[2],M[3],M[4],M[5],M[6],M[7],M[8],M[9],M[10],M[11],M[12],M[13],M[14],M[15],M[0],M[1]},S,SHO[2]);
mux16to1 T4({M[3],M[4],M[5],M[6],M[7],M[8],M[9],M[10],M[11],M[12],M[13],M[14],M[15],M[0],M[1],M[2]},S,SHO[3]);
mux16to1 T5({M[4],M[5],M[6],M[7],M[8],M[9],M[10],M[11],M[12],M[13],M[14],M[15],M[0],M[1],M[2],M[3]},S,SHO[4]);
mux16to1 T6({M[5],M[6],M[7],M[8],M[9],M[10],M[11],M[12],M[13],M[14],M[15],M[0],M[1],M[2],M[3],M[4]},S,SHO[5]);
mux16to1 T7({M[6],M[7],M[8],M[9],M[10],M[11],M[12],M[13],M[14],M[15],M[0],M[1],M[2],M[3],M[4],M[5]},S,SHO[6]);
mux16to1 T8({M[7],M[8],M[9],M[10],M[11],M[12],M[13],M[14],M[15],M[0],M[1],M[2],M[3],M[4],M[5],M[6]},S,SHO[7]);
mux16to1 T9({M[8],M[9],M[10],M[11],M[12],M[13],M[14],M[15],M[0],M[1],M[2],M[3],M[4],M[5],M[6],M[7]},S,SHO[8]);
mux16to1 T10({M[9],M[10],M[11],M[12],M[13],M[14],M[15],M[0],M[1],M[2],M[3],M[4],M[5],M[6],M[7],M[8]},S,SHO[9]);
mux16to1 T11({M[10],M[11],M[12],M[13],M[14],M[15],M[0],M[1],M[2],M[3],M[4],M[5],M[6],M[7],M[8],M[9]},S,SHO[10]);
mux16to1 T12({M[11],M[12],M[13],M[14],M[15],M[0],M[1],M[2],M[3],M[4],M[5],M[6],M[7],M[8],M[9],M[10]},S,SHO[11]);
mux16to1 T13({M[12],M[13],M[14],M[15],M[0],M[1],M[2],M[3],M[4],M[5],M[6],M[7],M[8],M[9],M[10],M[11]},S,SHO[12]);
mux16to1 T14({M[13],M[14],M[15],M[0],M[1],M[2],M[3],M[4],M[5],M[6],M[7],M[8],M[9],M[10],M[11],M[12]},S,SHO[13]);
mux16to1 T15({M[14],M[15],M[0],M[1],M[2],M[3],M[4],M[5],M[6],M[7],M[8],M[9],M[10],M[11],M[12],M[13]},S,SHO[14]);
mux16to1 T16({M[15],M[0],M[1],M[2],M[3],M[4],M[5],M[6],M[7],M[8],M[9],M[10],M[11],M[12],M[13],M[14]},S,SHO[15]);
endmodule
