`timescale 1ns/1ns
module barrel16tb();
logic [15:0]m=16'b0100100100100100;
logic [3:0]ss=4'b0000;
wire sho[15:0];
barrel16 UUT(m,ss,sho);
initial begin
#150 ss=4'b0010;
#150 ss=4'b0110;
#150 ss=4'b0100;
#150 ss=4'b1100;
#150 ss=4'b1110;
#150 ss=4'b1111;
#150 ss=4'b1011;
#150 m=16'b0100100101100100;
#150 m=16'b0100110101100100;
#150 m=16'b0100100100100100;
#150 m=16'b0100100100100110;
#150 m=16'b0100100110100100;
#150 m=16'b0110100100100100;
#150 ss=4'b1010;
#150 ss=4'b0010;
#150 $stop;
end
endmodule 